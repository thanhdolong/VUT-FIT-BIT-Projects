Nahradte obsahem souboru cpu.vhd nachazejiciho se v adresari fpga
